module pc (
	
	input wire CLK;

	);
